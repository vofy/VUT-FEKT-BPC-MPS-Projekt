BPC-MPS – Projekt

Vinp vin_p 0 DC 15
Vinn 0 vin_n DC 15

Xref        vin_p       0           ref_trim ref_vout REF-02/AD
Xout_adj    ref_vout    ref_trim    0                 OUT_ADJ
Rref_vout   ref_vout    opamp_inv                     50k
Xopamp      div_high    opamp_inv   vin_p  vin_n vout OP-97/LT
Rfeedback   opamp_inv   vout                          50k
Rdiv_vout   ref_vout    div_high                      12.5k
Rpot        div_high    div_low                       25k
Rdiv_gnd    div_low     0                             12.5k

.DC Vinp 0 60V .5V
.PROBE V([vout])

.LIB "lib/anlg_dev.lib"
.LIB "lib/linear_tech.lib"
.LIB "lib/subckts.lib"

.END